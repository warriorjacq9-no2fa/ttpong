module sprite #(

)
(
    input reg [10:0] x, y,
    output wire [3:0] r, g, b,
    output wire en
);

    assign en = ()

endmodule